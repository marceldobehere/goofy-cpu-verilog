module GoofyCore (

);

endmodule